library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity registro1 is
	Port(
		reloj : in STD_LOGIC;
		edo_sig : in std_logic_vector (2 downto 0);  --Liga
		entrada : in std_logic_vector ( 2 downto 0); --Los switch
		direccion : out std_logic_vector (5 downto 0));
end registro1;


architecture Behavioral of registro1 is
	begin
		process(reloj)
		begin
			if(rising_edge(reloj)) then
				direccion <= edo_sig & entrada;
			end if;
		end process;
end Behavioral;